----------------------------------------------------------------------------------
-- Project Name: Ping Pong Game
-- Brief: This module is the one that does the painting job. It contains the dynamic
--        position data belonging to different objects, it scans the screen and compares
--        the positions of the cursors with the position data, then it colors the screen
--        in the desired intersections. 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.Constants.all;

entity Sync is
  Port (clock, left, right, start: in std_logic;     
        difficultyControl: in std_logic_vector(1 downto 0);  
        hSync, vSync: out std_logic;
        r, g, b: out std_logic_vector(3 downto 0));        
end Sync;

architecture Behavioral of Sync is
--Defitions of the bitmaps for different images, they will be stored in the ROM 
type BITMAP1 is array (0 to 60) of std_logic_vector(0 to 299);
type BITMAP2 is array (0 to 46) of std_logic_vector(0 to 399);
type BITMAP3 is array (0 to 164) of std_logic_vector(0 to 199);
type BITMAP4 is array (0 to 63) of std_logic_vector(0 to 399);
--Synchronization Signals
signal hPosCurrent, hPosNext: integer range 1 to TOT_H;
signal vPosCurrent, vPosNext: integer range 1 to TOT_V;
--RGB Signals
signal rgbCurrent, rgbNext: std_logic_vector(11 downto 0);
--Intermediate Signals 
signal messageVisible, paddleVisible, ballVisible, frameVisible, paddleAIVisible, result1Visible, result2Visible, logoVisible, gameLabelVisible, borderVisible: boolean;
signal paddleCursor, paddleAICursor: integer range (FP_H + SP_H + BP_H + 1) to (TOT_H - PADDLE_WIDTH):= FP_H + SP_H + BP_H + VIS_H / 2 - (PADDLE_WIDTH + 1) / 2;
signal paddleLeft, paddleRight, paddleAILeft, paddleAIRight: integer range 0 to PRESCALER_PADDLE:= 0;
signal ballCursorX: integer range (FP_H + SP_H + BP_H + 1) to (TOT_H - BALL_SIDE);
signal ballCursorY: integer range (FP_V + SP_V + BP_V + 1) to (TOT_V - BALL_SIDE);
signal ballMovementCounter: integer:= 0;
signal ballMovement: std_logic:= '0';
signal playing: std_logic;
signal newGame, AIWins, playerWins: std_logic;
signal result1, result2: BITMAP1;
signal message: BITMAP2;
signal logo: BITMAP3;
signal gameLabel: BITMAP4;
signal paddleWidth: integer:= PADDLE_WIDTH; 
--Component that provides information about the balls position and game logic
component BallController is
    Port (start, move: in std_logic;
          paddleWidth: in integer;
          paddlePos, paddleAIPos: in integer range TOT_H - VIS_H + 1 to TOT_H - PADDLE_WIDTH;
          xPos: out integer range TOT_H - VIS_H + 1 to TOT_H - BALL_SIDE;
          yPos: out integer range TOT_V - VIS_V + 1 to TOT_V;
          newGame, play, AIWon, playerWon: out std_logic);
end component;
begin
    ballControl: BallController 
        port map (start => start,
                  move => ballMovement, 
                  paddleWidth => paddleWidth,
                  paddlePos => paddleCursor, 
                  paddleAIPos => paddleAICursor,
                  xPos => ballCursorX,
                  yPos => ballCursorY,
                  newGame => newGame, 
                  play =>  playing,
                  AIWon => AIWins,
                  playerWon => playerWins);
    --Bitmap assignments for the images             
    result1 <= ("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011000011111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110000001111111",
                "111111111111111100000001111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000001111111000000000111111100000000011111111111111111111001111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111110011001000000111111",
                "111111111111100000111000001111111111111111111111111111111000010000011111111111111111111111111111111111111111111111110000100000111111000010000011111100001000001111111111111100000000000111111111111111111111111000001110000011111111111111111111111111111111111111111111111111111111111100110111000000111111",
                "111111111110001111000111100111111111111111111111111111111010010110001111111111111111111111111111111111111111111111110110100100011111011010010001111101001011000111111111111000111111110001111111111111111111110011111001111000111111111111111111111111111111111111111111111111111111111001101100000000111111",
                "111111111100111000000000110001111111111111111111111111111010010110000111111111111111111111111111111111111111111111110110100100001111011010010000111101001011000011111111100011100000001110011111111111111111000110000000001110011111111111111111111111111111111111111111111111111111111011011001000000111111",
                "111111111001100011111110001100111111111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111111001110011111100011001111111111111110011000111111100011001111111111111111111111111111111111111111111111111111110010010011000000111111",
                "111111110011001110000011100110011111111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111110011001110000111001100111111111111100110011100000011001100111111111111111111111111111111111111111111111111111110110100100000000111111",
                "111111110110011000111000110011011111111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111110110010000000000110010011111111111101100110001110000100110011111111111111111111111111111111111111111111111111100100101100000000111111",
                "111111100100100111111111001001001111111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111101100100011111110011011001111111111001001100111111110010011001111111111111111111111111111111111111111111111111100101101000000000111111",
                "111111001001001100000001101101100111111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111001001001100000011001101100111111111011011011000000011001001000111111111111111111111111111111111111111111111111100101001000000000111111",
                "111111001011011000000000110110100011111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111011011011000000000100100100011111110010010010000000001101101100011111111111111111111111111111111111111111111111101101001000000001111111",
                "111111011010010000000000010010110001111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001111010010010000000000010110100001111110110100100000000000100100100011111111111111111111111111111111111111111111111101101001000000011111111",
                "111111010010100000000000011010010000111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010010100000000000010010110001111110100100100000000000010100100001111111111111111111111111111111111111111111111101101001000000111111111",
                "111110010110100000000000001010010000111111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010110100000000000011010010000111110100101000000000000010110100000111111111111111111111111111111111111111111111101101001000000111111111",
                "111110010110100000000011001011010000011111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000000000001010010000011110100101000000000110010010100000111111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000001111001011010000011111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000001111001010010000011110100101000000011111010010100000111111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000011111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000011111001010010000011110100101000000011111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000011111001010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000011111001010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000011111001010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000000000001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110111111111111111011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110111111111111111011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110000000000000000011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111000011111111101101001000001111111111",
                "111110010111111111111111111111010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111100011001111111101101001000001111111111",
                "111110010110000000000000000011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111101111100111111101101001000001111111111",
                "111110010110111111111111111011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111001000110011111101101001000001111111111",
                "111110010110110000000000011011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111011010010001111101101001000001111111111",
                "111110010110100000000000001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111001000110000111101101001000001111111111",
                "111110010110100000000000001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111001101100000011101101001000001111111111",
                "111110010110100000000000001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111100111000000011101101001000001111111111",
                "111110010110100000000000001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111110000000000011101101001000001111111111",
                "111110010110100000000000001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111000000000011101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111100000000011101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111110000000011101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000111011010010000011101001011000001110010100100000111111001010010000011110100101000000111111010010100000011111111111111111111111111111111111000000111101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110110100100000110010011010000011101001011000001110010010100000111111010010010000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110010100100000110110111011000011001001010000001111010010010000111110010010110000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000001111111111111111111010010110000011111111111111111111111111111111111111111111110010110110000000100111001000010011011010000001111011011011000111100100100100000011110100101000000111111010010100000011111111111111111111111111111111111111111111101101001000001111111111",
                "111110010110100000011111001011010000001111100001111111111010010110000011111100001111111111111111111111111111111111111010010011000001001101100100000110010010000001111001001001100000001101101100000011110100101000000111111010010100000011111111111111111111111111111110000011111111100101001000001111111111",
                "111110010110100000011111001011010000001111001100111111111010010110000011110001100111111111111111111111111111111111111011011001111110011000110011111100110110000001111101100100111000110001001000000011110100101000000111111010010100000011111111111111111111111111111100111001111111100101001000001111111111",
                "111110010110100000011111001011010000001110011110011111111010010110000011110111110011111111111111111111111111111111111001001100001000110000011000100001100100000001111100110010001111100110011000000011110100101000000111111010010100000011111111111111111111111111111101111100111111100101101000001111111111",
                "111110010110100000011111001011010000001110100001001111111010010110000011100100001001111111111111111111111111111111111100100111000001100111001110000111001000000001111110011001100000001100110000000011110100101000000111111010010100000011111111111111111111111111111001000110011111110100100100001111111111",
                "111110010110100000011111001011010000001110101101000111111010010110000011100101001000111111111111111111111111111111111110110001111110001101100011111100011000000001111111001100111111111001100000000011110100101000000111111010010100000011111111111111111111111111111011010010001111110010110010001111111111",
                "111110010110100000011111001011010000001110100001000011111010010110000011100100011000011111111111111111111111111111111110001100000000011000110000000001100000000011111111100110000000000111000000000111110100101000000111111010010100000011111111111111111111111111111001000110000111110010011001000111111111",
                "111110010110100000011111001011010000001110011110000001111010010110000011110111110000001111111111111111111111111111111111100111111111100000001111111111000000000011111111110011110000011100000000000111110100101000000111111010010100000011111111111111111111111111111101111100000011111001001100000111111111",
                "111110010000100000011111001000010000001111000000000000111010010000000011110000000000001111111111111111111111111111111111110000011100000000000001110000000000000011111111111000011111110000000000001111110100101000000111111010010100000011111111111111111111111111111100000000000011111101100110000011111111",
                "111110000000000000011111000000000000001111100000000000111000000000000011111100000000000111111111111111111111111111111111111000000000000000000000000000000000000111111111111100000000000000000000011111110000000000000111111000000000000011111111111111111111111111111110000000000011111100110001000001111111",
                "111111000000000000011111100000000000001111110000000000111100000000000011111110000000000111111111111111111111111111111111111100000000000000000000000000000000001111111111111110000000000000000000111111111000000000000111111100000000000011111111111111111111111111111111000000000011111110001100000000111111",
                "111111100000000000011111110000000000001111111000000000111110000000000011111111000000001111111111111111111111111111111111111110000000000000000100000000000000011111111111111111000000000000000001111111111100000000000111111110000000000011111111111111111111111111111111100000000011111111100111000000111111",
                "111111110000000000011111111000000000001111111100000001111111000000000011111111100000001111111111111111111111111111111111111111000000000000011110000000000000111111111111111111100000000000000011111111111110000000000111111111000000000011111111111111111111111111111111110000000011111111110001000000111111",
                "111111111000000000011111111100000000001111111110000011111111100000000011111111110000011111111111111111111111111111111111111111110000000001111111100000000111111111111111111111111000000000001111111111111111000000000111111111100000000011111111111111111111111111111111111100001111111111111000000000111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");          
    result2 <= ("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011001111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011001111111111111",
                "111100000000011111111100000000011111111111111000000000111111111111111000000000111111111000000000111111111111111111111111111111100000000011111100000000011111100000000011111111111111100000000011111111111111111111111000000000001111111111111111111111111111111111111111111111111111111011001100111111111111",
                "111101101010001111111101001010001111111111100011111110001111111111111001010110011111111011010100011111111111111111111111111111101101010001111101101011001111101001010001111111111110001111111000111111111111111111110011111111100011111111111111111111111111111111111111111111111111111000110110111111111111",
                "111101101010000111111101001010000111111110011110000011100111111111111001010110001111111011010100001111111111111111111111111111101101010000111101101011000111101001010000111111111001110000001110011111111111111111001110000000011001111111111111111111111111111111111111111111111111111010011010011111111111",
                "111101101010000011111101001010000011111100110001111100011001111111111001010110000111111011010100000111111111111111111111111111101101010000011101101011000011101001010000011111110011000111110001100111111111111110011001111111000100111111111111111111111111111111111111111111111111111001001001001111111111",
                "111101101010000001111101001010000011111001100111000111001100111111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011111100110011100011100110011111111111100110111000001110010011111111111111111111111111111111111111111111111111000100101000111111111",
                "111101101010000001111101001010000011111011011000000000110110111111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011111101101100000000011011011111111111101101100011100011001001111111111111111111111111111111111111111111111111100110100100011111111",
                "111101101010000001111101001010000011110110110011111110011011011111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011111011011001111111001101101111111111011011001110111100100100111111111111111111111111111111111111111111111111110010100100001111111",
                "111101101010000001111101001010000011100100100100000001001001001111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110010010010000000100100100111111111010010010000000110110110011111111111111111111111111111111111111111111111111010010100001111111",
                "111101101010000001111101001010000011101101001000000000100101100111111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110110100100000000010010110011111110010100100000000011010010001111111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011101001010000000000010100100011111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110100101000000000001010010001111110100101000000000001001010000111111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011101010010000000000010010100001111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011110101001000000000001001010000111110100101000000000001001010000111111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000000000011010100000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101001000000000001101010000111110101001000000000000101011000011111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000000111011010100000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101001000000011101101010000011110101001000000011100101011000011111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000001111011010110000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000000111101101010000011110101001000000111100101011000011111111111111111111111111111111111111111111111010010100000111111",
                "111101101010000001111101001010000011001010010000011111011010110000111001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000011110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111100101011000001111101001010000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111100101001000001111101010010000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111110101101000001111001010010000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111110100100100001110010010100000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111110010110011000000100100100000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111111011011001111111001001000000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111110001111111111111010010100000111111",
                "111111001001110000000010011000000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111000100011111111111010010100000111111",
                "111111100100011110111100110000000011001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111011111011111111111010010100000111111",
                "111111110011000111100001100000000111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111110010001001111111111010010100000111111",
                "111111111001110001000110000000000111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111110110101000111111111010010100000111111",
                "111111111100001101011000000000001111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111110010001000011111111010010100000111111",
                "111111111110001101010000000000001111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111011111000001111111010010100000111111",
                "111111111111001101010000000000011111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111000100000000111111010010100000111111",
                "111111111111101101010000000000111111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111100000000000111111010010100000111111",
                "111111111111101101010000000011111111001010010000011111011010110000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111000000000111111010010100000111111",
                "111111111111101101010000001111111111001010010000011111011010100000011001010110000011111011010100000011111111111111111111111111101101010000001101101011000001101001010000011100101011000001111101101010000001110101001000001111100101011000001111111111111111111111111111111100000001111111010010100000111111",
                "111111111111101101010000001111111111001010010000011111011010100000011001010010000011111010010100000011111111111111111111111111101101010000001101101011000001101001010000011100101001000001111101101010000001110101001000001111100101011000001111111111111111111111111111111110000001111111010010100000111111",
                "111111111111101101010000001111111111101010010000011111010010100000011001010010000011111010010100000011111111111111111111111111101101010000001101001001000001101001010000011110101001000001111101001010000001110101001000001111100101011000001111111111111111111111111111111111000111111111010010100000111111",
                "111111111111101101010000001111111111101001010000011111010110100000011101011010000011110010100100000011111111111111111111111111100101001000001001011101000001101001010000011110100101000001111101011010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111111111111101101010000001111111111101101001000011110010100100000011101101001000011100100100100000011111111111111111111111111100101001000000011011101100001001011010000011110110100100001111001010010000001110101001000001111100101011000001111111111111111111111111111111111111111111111010010100000111111",
                "111111111111101101010000001111111111100100101100010000101101100000011100101101100000001101101000000011111111111111111111111111110100100100000110110110100000010010010000011110010010110001000010110100000001110101001000001111100101011000001111111111111111111111111111110001111111111111010010100000111111",
                "111111111111101101010000001111111111110110110111000011001001000000011110110110011111111001001000000111111111111111111111111111110100110011111100100010011111100110100000011111011010011100001100100100000001110101001000001111100101011000001111111111111111111111111111000100011111111111010110100000111111",
                "111111111111101101010000001111111111110010011001111100110010000000111110010011000111000110010000000111111111111111111111111111110010011000110001100011000110001100100000011111001001100111110011001000000011110101001000001111100101011000001111111111111111111111111111011111011111111110010100100000111111",
                "111111111111101101010000001111111111111001001100000001100110000000111111001001110000011100100000000111111111111111111111111111111011001110000110011101110000111001000000011111100100110000000110011000000011110101001000001111100101011000001111111111111111111111111110010001001111111100100101000000111111",
                "111111111111101101010000001111111111111100100011111111001100000000111111100110011111110001000000000111111111111111111111111111111101100011111100110100011111100010000000011111110010001111111100110000000011110101001000001111100101011000001111111111111111111111111110110101000111111001001001000000111111",
                "111111111111101101010000001111111111111110011000000000110000000000111111110011000000000110000000001111111111111111111111111111111100111000000001100011000000001100000000011111111001100000000011000000000111110101001000001111100101011000001111111111111111111111111110010001000011111010011011000000111111",
                "111111111111101101010000001111111111111111001111000111100000000001111111111000111111111000000000001111111111111111111111111111111111001111111110000000111111111000000000111111111100111100011110000000000111110101001000001111100101011000001111111111111111111111111111011110000001111000110110000000111111",
                "111111111111100001000000001111111111111111100001111100000000000011111111111100000000000000000000011111111111111111111111111111111111100000000000000000000000000000000000111111111110000111110000000000001111110100000000001111100001000000001111111111111111111111111111000000000000111011101100000000111111",
                "111111111111100000000000001111111111111111110000000000000000000011111111111110000000000000000000111111111111111111111111111111111111110000000000000000000000000000000001111111111111000000000000000000011111110000000000001111110000000000001111111111111111111111111111110000000000111010011000000001111111",
                "111111111111110000000000001111111111111111111000000000000000000111111111111111000000000000000001111111111111111111111111111111111111111000000000000000000000000000000011111111111111100000000000000000011111111000000000001111111000000000001111111111111111111111111111111000000000111001110000000001111111",
                "111111111111111000000000001111111111111111111100000000000000011111111111111111100000000000000011111111111111111111111111111111111111111100000000000000110000000000000111111111111111110000000000000001111111111100000000001111111100000000001111111111111111111111111111111100000001111011000000000011111111",
                "111111111111111100000000001111111111111111111111000000000000111111111111111111111000000000001111111111111111111111111111111111111111111110000000000011111000000000001111111111111111111100000000000011111111111110000000001111111110000000001111111111111111111111111111111110000001111000000000000011111111",
                "111111111111111111000000011111111111111111111111110000000111111111111111111111111111000001111111111111111111111111111111111111111111111111110000011111111111000001111111111111111111111111000000011111111111111111000000001111111111000000001111111111111111111111111111111111000111111000000000000111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000001111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");          
	message <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111000000001111111111111111111111100000000111111111111111000000001111110000000001111100000000111111111111111111111111111111111111110000000011111111111111111111111000000001111111111111111111111000000001111110000000001111111111111111111100000000011111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111110000000011111111111111111111111111111111",
                "1111111111100111111110001111111111111111100011111111001111111111111010110100111110100101000111101011010011111111111111111111111111111111111001111111000111111111111111111100111111110011111111111111111100111111100011000111111100111111111111111110001111111100111111111111111111111111111111111111111111111111111011111111111111100111111111111111111111111111111111001111111000111111111111111111111111111111",
                "1111111110011100000001100111111111111111001100000000110011111111111010110100011110100101000011101011010001111111111111111111111111111111100111000000110001111111111111110011100000001100111111111111110011000000001000011000000011001111111111111100110000000011001111111111111111111111111111111111111111111111111010000000000000011001111111111111111111111111111100111000000110011111111111111111111111111111",
                "1111111100110011111100010011111111111110011001111110011001111111111010110100001110100101000001101011010000111111111111111111111111111111001100011110001100111111111111100110011111100010011111111111110100011111100100100111111000100111111111111001100111111001100111111111111111111111111111111111111111111111111010111111111111001100111111111111111111111111111001100011110001101111111111111111111111111111",
                "1111111001001110000011001001111111111100100110000001100100111111111010110100000110100101000001101011010000011111111111111111111111111110010011100001100110011111111111001001110000011001001111111111101001110000110011001100001110010011111111110010011000000110010011111111111111111111111111111111111111111111111010100000000000110010011111111111111111111111110010011100001110110111111111111111111111111111",
                "1111111010011001111000100100111111111001001100111100110010011111111010110100000110100101000001101011010000011111111111111111111111111110100110001100011011011111111111010011001111000100100111111111001011000110001000010001110011001001111111100100110011110011001001111111111111111111111111111111111111111111111010101111111110011001011111111111111111111111110100110001100011011011111111111111111111111111",
                "1111110110100110000110010010011111111011010011100111001011001111111010110100000110100101000001101011010000011111111111111111111111111101101001111111101101001111111110110100110001110010010011111111010010011001100100100110001001101000111111101101001110011100101100111111111111111111111111111111111111111111111010101100000001100101101111111111111111111111101101001111111101101001111111111111111111111111",
                "1111110101101000000001001010001111110010110110000001101101000111111010110100000110100101000001101011010000011111111111111111111111111001011011000000110100100111111110101101000000001001010001111111010100100000010111101000000100101000111111001011011000000110110100011111111111111111111111111111111111111111111010101000000000010110100111111111111111111111001011011000000110110100111111111111111111111111",
                "1111100101010000000000101001000111110110101100000000110100100011111010110100000110100101000001101011010000011111111111111111111111111011010110000000011010100011111101101010000000000101001000111110010101000000010011001000000010100100011111011010110000000011010010001111111111111111111111111111111111111111111010101000000000001010100011111111111111111111010010110000000011010100011111111111111111111111",
                "1111101001010000000000100101000111110101101000000000010010100011111010110100000110100101000001101011010000011111111111111111111111111010110100000000001010010001111101001010000000000100101000111110100101000000001011010000000010010100001111010110100000000001001010001111111111111111111111111111111111111111111010101000000000001010010001111111111111111111010110100000000001011010001111111111111111111111",
                "1111101010010000000000010101000011110101001000000000011010100001111010110100000110100101000001101011010000011111111111111111111111111010100100000000001001010000111101010010000000000010101000011110100101000000001011010000000010010100001111010101100000000001101010000111111111111111111111111111111111111111111010101000000000001101010000111111111111111111010100100000000001001010000111111111111111111111",
                "1111101010010000000010010101000011110101010000000001011010100001111010110100000110100101000001101011010000011111111111111111111111111010101000000000101101010000111101010110000000010010101000011110100101000000001011010000000010010100001111010101000000000101101010000111111111111111111111111111111111111111111010101000001111101101010000111111111111111111010101000000000101101010000111111111111111111111",
                "1111101010110000001110010101000001110101010000000111000000000000111010110100000110100101000001101011010000011111111111111111111111111010101000000011100000000000011101010110000001110010101000001110100101000001101011010000001010010100000111010101000000011100000000000011111111111111111111111111111111111111111010101000001111101101010000111111111111111111010101000000011100000000000111111111111111111111",
                "1111101010110000011110010101000001110101010000001111100000000000111010110100000110100101000001101011010000011111111111111111111111111010101000000111110000000000011101010110000011110010101000001110100101000001101011010000011010010100000111010101000000111110000000000011111111111111111111111111111111111111111010101000001111101101010000011111111111111111010101000000111110000000000011111111111111111111",
                "1111101010110000011110010101000001110101010000001111110000000000111010110100000110100101000001101011010000011111111111111111111111111010101000000111111000000000011101010110000011110010101000001110100101000001101011010000011010010100000111010101000000111111000000000011111111111111111111111111111111111111111010101000001111101001010000011111111111111111010101000001111111000000000011111111111111111111",
                "1111101010110000111110010101000001110101010000011111111000000000111010110100000110100101000001101011010000011111111111111111111111111010101000001111111100000000011101010110000111110010101000001110100101000001101011010000011010010100000111010101000001111111100000000011111111111111111111111111111111111111111010101000001111011010010000011111111111111111010101000001111111100000000011111111111111111111",
                "1111101010110000111110010101000001110101010000001111111100000000111010110100000110100101000001101011010000011111111111111111111111111010101000000111111100000000011101010110000011110010101000001110100101000001101011010000011010010100000111010101000000111111110000000011111111111111111111111111111111111111111010101000000000010010100000011111111111111111010101000001111111110000000011111111111111111111",
                "1111101010110000111110010101000001110101011000000000001111111111111010110100000110100101000001101011010000011111111111111111111111111010101000000000000000000011111101010110000000000110101000001110100101000001101011010000011010010100000111010101100000000000111111111111111111111111111111111111111111111111111010101100000011100100100000011111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101011111111111000111111111111010110100000110100101000001101011010000011111111111111111111111111010101000000111111111110001111101010011111111111110101000001110100101000001101011010000011010010100000111010101111111111100011111111111111111111111111111111111111111111111111010101111111110001101000000011111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101000000000000000011111111111010110100000110100101000001101011010000011111111111111111111111111010101000000000000000010000111101010000000000000000101000001110100101000001101011010000011010010100000111010100000000000000001111111111111000111111111111111111111111111111111010100000000000011011000000011111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101111111111111000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000000111111111010000011101011111111111111111101000001110100101000001101011010000011010010100000111010111111111111100000111111111110011001111111111111111111111111111111010111111111111110010000000111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101000000000000000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000000000000001010000011101010000000000000000101000001110100101000001101011010000011010010100000111010100000000000000000111111111101111100111111111111111111111111111111010100000000000111001000000111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101011111111111000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000000111111001010000011101010111111111111110101000001110100101000001101011010000011010010100000111010101111111111100000111111111101000100011111111111111111111111111111010101111111110001100100000111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101011000000000000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000000000001101010000011101010110000000000010101000001110100101000001101011010000011010010100000111010101100000000000000111111111101010100001111111111111111111111111111010101100000001100100100001111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101010000000000000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000000000000101010000011101010110000000000010101000001110100101000001101011010000011010010100000111010101000000000000000111111111101000100001111111111111111111111111111010101000000000110010000001111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101010000000000000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000001000000101010000011101010110000000000010101000001110100101000001101011010000011010010100000111010101000000000000000111111111100111000000111111111111111111111111111010101000000000011010010001111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101010000000000000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000001100000101010000011101010110000000000010101000001110100101000001101011010000011010010100000111010101000000000000000111111111110000000000111111111111111111111111111010101000000000001011010000111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101010000000000000001111111111010110100000110100101000001101011010000011111111111111111111111111010101000001110000101010000011101010110000000000010101000001110100101000001101011010000011010010100000111010101000000000000000111111111111000000000011111111111111111111111111010101000000000001101010000111111111111111111010101000001111111111111111111111111111111111111",
                "1111101010110000111110010101000001110101010000011111000000000111111010110100000110100101000001101011010000011111111111111111111111111010101000001111100101010000011101010110000111110010101000001110100101000001101011010000011010010100000111010101000001111100000000011111111100000000111111111111111111111111111010101000001111101101010000011111111111111111010101000001111100000000011111111111111111111111",
                "1111101010110000111110010101000001110101010000011111011010100011111010110100000110100101000001101011010000011111111111111111111111111010101000001111101101010000011101010110000111110010101000001110100101000001101011010000011010010100000111010101000001111101101010001111111110000000111111111111111111111111111010101000001111101101010000011111111111111111010101000001111101101010001111111111111111111111",
                "1111101010110000111110010101000001110101001000011111011010100001111010110100000110101101000001101011010000011111111111111111111111111010100100001111101001010000011101010110000111110010101000001110100101000001101011010000011010010100000111010100100001111101101010000111111111100001111111111111111111111111111010101000001111101101010000011111111111111111010101000001111101001010000111111111111111111111",
                "1111101010110000111110010101000001110101101000011110010010100000111010010100000100101101000001101010010000011111111111111111111111111010110100001111101001010000011101010110000111110010101000001110100101000001101011010000011010010100000111010110100001111001001010000011111111111111111111111111111111111111111010101000001111101011010000011111111111111111010100100001111101001010000011111111111111111111",
                "1111101010110000111110010101000001110110101000011100110100100000111010010100000001001100100001001010010000011111111111111111111111111010010100001111001010110000011101010110000111110010101000001110100101000001101011010000011010010100000111011010100001110011010110000011111111111111111111111111111111111111111010101000001111011010100000011111111111111111010010100001111011010000000011111111111111111111",
                "1111101010110000111110010101000001110010110110000001100101000000111001010010000011011010010000010010100000011111111111111111111111111001011010000100010010100000011101010110000111110010101000001110100101000001101011010000011010010100000111001011011000000110010100000011111000111111111111111111111111111111111010101000000000110110100000011111000111111111001011010000000110110100000011111000111111111111",
                "1111101010110000111110010101000001111011011001111111001011000000111101001001111110110011001111100100100000011111111111111111111111111101101001110001100100100000011101010110000111110010101000001110100101000001101011010000011010010100000111101101000111111100101100000011110010001111111111111111111111111111111010101111111111101101100000011110010011111111101101001100011100100100000011110010001111111111",
                "1111101010110000111110010101000001111101001100001000110010000000111100101100000001100001100000001101100000011111111111111111111111111110100110011110001001000000011101010110000111110010101000001110100101000001101011010000011010010100000111110100110000100011001000000011100111101111111111111111111111111111111010100111111100011011000000011101111101111111100100110011110001001000000011100111101111111111",
                "1111101010110000111110010101000001111100100111100011100100000000111110100011100111001100111000110001000000111111111111111111111111111110010011000000110010000000011101010110000111110010101000001110100101000001101011010000011010010100000111110010011110001110110000000011101000100111111111111111111111111111111010100000000011110110000000111101000100111111110010011000000110010000000111101000100111111111",
                "1111101010110000111110010101000001111110011000111110011000000001111110011000111100010010001111000110000000111111111111111111111111111111001100111111000100000000111101010110000111110010101000001110100101000001101011010000011010010100000111111001100011111001100000000111101010100011111111111111111111111111111010111111111110001100000000111001010100011111111001100111111000100000000111101010100011111111",
                "1111101010110000111110010101000001111111001110000001110000000001111111001110000001100001100000011100000000111111111111111111111111111111100110000000011000000000111101010110000111110010101000001110100101000001101011010000011010010100000111111100111000000111000000000111101100100001111111111111111111111111111010000000000000111000000000111101000100001111111100110000000011000000000111101100100001111111",
                "1111101010110000111110010101000001111111100001111111000000000011111111110011111110000000011111110000000000111111111111111111111111111111110001111111100000000001111101010110000111110010101000001110100101000001101011010000011010010100000111111110000111111100000000001111100111000000111111111111111111111111111011111111111111000000000001111100111000000111111110001111111100000000001111100111000000111111",
                "1111100000000000111110000000000001111111110000000000000000000111111111111000000000000000000000000000000001111111111111111111111111111111111000000000000000000011111100000000000111110000000000001110000000000001100000000000011000000000000111111111000000000000000000011111110000000000111111111111111111111111111000000000000000000000000011111110000000000111111111000000000000000000011111110000000000111111",
                "1111100000000000111111000000000001111111111000000000000000000111111111111100000000000000000000000000000011111111111111111111111111111111111100000000000000000011111100000000000111111000000000001111000000000001110000000000011100000000000111111111100000000000000000111111111000000000011111111111111111111111111000000000000000000000000111111111000000000111111111100000000000000000111111111000000000011111",
                "1111110000000000111111100000000001111111111110000000000000011111111111111110000000000000000000000000000111111111111111111111111111111111111110000000000000000111111110000000000111111100000000001111100000000001111000000000011110000000000111111111111000000000000001111111111110000000111111111111111111111111111100000000000000000000001111111111100000000111111111110000000000000001111111111110000000111111",
                "1111111000000000111111110000000001111111111111000000000000111111111111111111000000000001111000000000001111111111111111111111111111111111111111100000000000011111111111000000000111111110000000001111110000000001111100000000011111000000000111111111111100000000000011111111111111000000111111111111111111111111111110000000000000000000011111111111110000001111111111111100000000000011111111111111000000111111",
                "1111111100000000111111111000000001111111111111111000000011111111111111111111110000000111111110000001111111111111111111111111111111111111111111111000000001111111111111100000000111111111000000001111111000000001111110000000011111100000000111111111111111100000011111111111111111100011111111111111111111111111111111000000000000000011111111111111111100011111111111111111000000001111111111111111100011111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");          
logo <= (    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111",
             "11111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111",
             "11111111111111111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000001111111111111111111111111111111",
             "11111111111111111111111111111110000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111",
             "11111111111111111111111111111000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111",
             "11111111111111111111111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111",
             "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
             "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
             "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
             "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
             "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
             "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111",
             "11111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
             "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
             "11111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
             "11111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111100000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111110000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111000000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111100000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
             "11111111111110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111110000000000000000000000000000000000000000000000000000000000000000000001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
             "11111111111111000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
             "11111111111111100000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
             "11111111111111110000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
             "11111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
             "11111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
             "11111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
             "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
             "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
             "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
             "11111111111111111111000000000000000000000000000000000000000000000000000000000000000000011111001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
             "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111100011111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
             "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111100000111111110000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111",
             "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111100000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
             "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000011110000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
             "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011110000000001111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
             "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000011110000000000011111111000000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
             "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000111111000000000001111111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
             "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111111000000000000011111111000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
             "11111111111111111111111111100000000000000000000000000000000000000000000000000000000001111111111000000000000000111111110000000000000000000000000000000000000000000000000000000001111111111111111111111111",
             "11111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111111111111",
             "11111111111111111111111111111000000000000000000000000000000000000000000000000000001111111100111000000000000000000111111111000000000000000000000000000000000000000000000000000011111111111111111111111111",
             "11111111111111111111111111111100000000000000000000000000000000000000000000000000111111110001111000000000000000000001111111100000000000000000000000000000000000000000000000000111111111111111111111111111",
             "11111111111111111111111111111110000000000000000000000000000000000000000000000011111111000001111000000000000000000000111111111000000000000000000000000000000000000000000000001111111111111111111111111111",
             "11111111111111111111111111111111000000000000000000000000000000000000000000000111111110000001111000000000000000000000001111111110000000000000000000000000000000000000000000011111111111111111111111111111",
             "11111111111111111111111111111111100000000000000000000000000000000000000000011111111000000001111000000000000000000000000011111111000000000000000000000000000000000000000000111111111111111111111111111111",
             "11111111111111111111111111111111110000000000000000000000000000000000000001111111100000000001110000000000000000000000000001111111110000000000000000000000000000000000000001111111111111111111111111111111",
             "11111111111111111111111111111111111000000000000000000000000000000000000011111110000000000011110000000000000000000000000000011111111100000000000000000000000000000000000111111111111111111111111111111111",
             "11111111111111111111111111111111111100000000000000000000000000000000001111111100000000000011110000000000000000000000000000000111111110000000000000000000000000000000001111111111111111111111111111111111",
             "11111111111111111111111111111111111111000000000000000000000000000000111111110000000000000111110000000000000000000000000000000001111111100000000000000000000000000000011111111111111111111111111111111111",
             "11111111111111111111111111111111111111100000000000000000000000000011111111000000000000000111100000000000000000000000000000000000111111111000000000000000000000000001111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111000000000000000000000000111111110000000000000001111100000000000000000000000000000000000001111111100000000000000000000000111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111110000000000000000000011111111000000000000000001111000000000000000000000000000000000000000011111111000000000000000000011111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111000000000000000001111111100000000000000000011111000000000000000000000000000000000000000001111111110000000000000001111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111000000000000111111111000000000000000000011110000000000000000000000000000000000000000000011111111110000000001111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111000000111111111111111111000000000000111110000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111110000001111100000000000000000000000111110000001111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111100000011111100000000000000000000001111111000001111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100000000000000000000001111111000000111111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111000001111111110000000000000000000001111111100000011111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111110000001111111100000000000000000000001111111110000011111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000000000000000111111111000001111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000000000000000000111111111000000111111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111000001111111111000000000000000000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111110000001111111110000000000001100000000000001111111110000011111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000001110000000000001111111110000001111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111000000111111111100000000000011110000000000000111111111000000111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000000111111000000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111110000001111111110000000000000111111100000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000001111111100000000000001111111110000001111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111100000011111111100000000000001111111110000000000000111111111000000111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111000000111111111000000000000011111111111000000000000111111111100000111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111110000001111111110000000000000111111111111000000000000011111111100000011111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111100000001111111110000000000000111111111111100000000000001111111110000001111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111100000001111111100000000000001111111111111110000000000000111111110000000111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111000000001111111000000000000011111111111111110000000000000111111110000000111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000000111110000000000000011111111111111111000000000000011111100000000011111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000000011100000000000000111111111111111111100000000000000110000000000001111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111100000000000000000000011111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111",
             "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

    gameLabel <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111000000000000000000000011111111111111111111111111111111000000011111111111111111111111111111111110000000000011111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111100000000001111111111111111111111111111111000000000011111111110000000000111111111111111111111111111111100000000000111111111111111111111111",
                  "1111111011111111111111111100000111111111111111111111111110000000000000011111111111111111111111111111000001111100000111111111111111111111111111100000111110000011111111111111111111111111111111111111111111111111111111111100000111100000011111111111111111111111111100000011111000001111111111111111111111111100000111110000111111000001111100000111111111111111111111111100000011111000001111111111111111111111",
                  "1111111011111111111111111111110001111111111111111111111000011111111110000111111111111111111111111100001111111111110001111111111111111111111110001111111111110000111111111111111111111111111111111111111111111111111111110001111111111110001111111111111111111111110000111111111111000111111111111111111111110001111111111110001100011111111111100011111111111111111111111000111111111111000011111111111111111111",
                  "1111111011000000000000000000011100111111111111111111110001111000000011110001111111111111111111111000111000000000011100111111111111111111111100011100000000111100011111111111111111111111111111111111111111111111111111000111100000000111100111111111111111111111100011100000000001110001111111111111111111100111000000000011100001110000000000111001111111111111111111100011100000000001110001111111111111111111",
                  "1111111011011111111111111110000110011111111111111111100111100000000000011000111111111111111111110011100001111110000110001111111111111111111001110000011100000110001111111111111111111111111111111111111111111111111110001110000111100001110001111111111111111111000110000111111000011100111111111111111111001100001111110000110011000011111100001100111111111111111111000110000111111000011100111111111111111111",
                  "1111111011011111111111111111100011001111111111111111001110011111111111001110011111111111111111100110001111111111100011000111111111111111110011000111111111100011000111111111111111111111111111111111111111111111111100011000111111111100011000111111111111111110011100111111111111001110011111111111111110011000111111111100011110001111111111000110011111111111111110011100011111111111001110011111111111111111",
                   "1111111011011000000000000000111001100111111111111110011100111000000011100011001111111111111111001100111100000000111001100111111111111111100110011110000000111001100011111111111111111111111111111111111111111111111000110011110000001111001100111111111111111100111001110000000011100011001111111111111110110001110000000111001100011000000001110011001111111111111100111001110000000011100011001111111111111111",
                  "1111111011011001111111111100001100110011111111111100111011100000000000111001100111111111111110011001110000111100001100110011111111111111001100111000000000001100110001111111111111111111111111111111111111111111111001100110000000000001100110011111111111111100110011000011110000110011000111111111111100100011000011100011100001110001111000111001100111111111111100110011000011110000111001100111111111111111",
                  "1111111011011011111111111111000110011001111111111100110010000111111110001100110011111111111110010011000111111111000110011001111111111110011001100011111111100110011000111111111111111111111111111111111111111111110011001100011111111000110011001111111111111001100110011111111110011001100011111111111101100110001111111001110001100111111110011100100011111111111001100110011111111110011101110011111111111111",
                  "1111111011011011000000000001110011001000111111111001100100011100000111000110110001111111111100110010001100000001110011001000111111111110010011000110000001110011001100011111111111111111111111111111111111111111110110011001110000001110011001000111111111110011001100110000000111001100110001111111111001001100110000001100110011001100000011001100110001111111111011001100111000000011001100110001111111111111",
                  "1111111011011011000000000000011001001100011111111001001100110000000001100010011000111111111100100110010000000000011001001100011111111100110010001100000000011001100100001111111111111111111111111111111111111111100110110011000000000011001001100011111111110010011001100000000001100110010000111111111001001100100000000110011010011000000001100110110000111111110011011001100000000001100110011000111111111111",
                  "1111111011011011000000000000001001100100001111110011001001100000000000010011001000011111111001101100100000000000001001100100001111111100100110010000000000001100100110000111111111111111111111111111111111111111101100100110000000000001101100100001111111110110010011000000000000110010011000011111111011001001100000000010011110010000000000100110010000011111110010011011000000000000110011011000011111111111",
                  "1111111011011011000000000000000100100100000111110010011001000000000000011001001000001111111001001101100000000000001100100110000111111101100100110000000000000110110010000111111111111111111111111111111111111111001101100100000000000000100100110000111111100110110010000000000000010011011000011111111011011001000000000011001110110000000000110010010000011111110110010010000000000000011011001000001111111111",
                  "1111111011011011000000000000000100110110000111110010010011000000000000001001101100001111111001001001000000000000000100110110000011111101101100100000000000000110010010000011111111111111111111111111111111111111001001101100000000000000110110010000011111100100110110000000000000011011001000001111110011011011000000000001001100100000000000010010010000001111100110110110000000000000011001001000001111111111",
                  "1111111011011011000000000000000110110110000011110110010010000000000000001101101100000111111011001001000000000000000110110010000011111001101100100000000000000010010010000001111111111111111111111111111111111111001001001100000000000000110010010000011111100100100100000000000000001001001000001111110011011011000000000001001100100000000000010010010000001111100100100110000000000000001001001100000111111111",
                  "1111111011011011000000000000000010110010000001110110110010000000000000001101100100000111111011011001000000000000000110110010000001111001001101100000000000000011011011000001111111111111111111111111111111111111001001001000000000000000010010010000001111100100100100000000000000001001001000000111110011011011000000000001101101100000000000010010011000000111100100100100000000000000001001101100000111111111",
                  "1111111011011011000000011111110010110010000001110110110010000000000111101101100100000011111011011001000000000111110110110010000001111001001101100000000001110010011011000000111111111111111111111111111111111111001001001000000000011110010010010000001111100100100100000000001111001001001000000111110011011011000000001101101101100000000010010010011000000111100100100100000000001111001001101100000011111111",
                  "1111111011011011000000011111110010110010000001110110110010000000011111101101100100000011111011011001000000001111110110110010000001111001001101100000000111110000000000000000111111111111111111111111111111111111001001001000000000111110000000000000000111100100100100000000011111001001001000000011110011011011000000011101101101100000000110010010011000000111100100100100000000011111000000000000000011111111",
                  "1111111011011011000000011111100110110110000001110110110010000000011111101101100100000011111011011001000000001111110110110010000000111001001101100000001111111000000000000000111111111111111111111111111111111111001001001000000001111110000000000000000111100100100100000000111111001001001000000011110011011011000000011101101101100000001110010010011000000111100100100100000000111111100000000000000011111111",
                  "1111111011011011000000011111100100110110000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111100000000000000111111111111111111111111111111111111001001001000000001111111100000000000000111100100100100000001111111001001001000000011110011011011000000011101101101100000001110010010011000000111100100100100000000111111110000000000000011111111",
                  "1111111011011011000000011111100100100110000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111110000000000000111111111111111111111111111111111111001001001000000011111111110000000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111111000000000000011111111",
                  "1111111011011011000000011111001001100100000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111111111000000000000111111111111111111111111111111111111001001001000000011111111111000000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111111100000000000001111111",
                  "1111111011011011000000011100011001101100000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111100000000000111111111111111111111111111111111111001001001000000011111111111000000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111111110000000000001111111",
                  "1111111011011011000000000001110011001000000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000000000000000111111111111111111111111111111111111001001001000000000000000000000000000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000011111000000000011111111",
                  "1111111011011011111111111111000110011000000000110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111111111000111111111111111111111111111111111111111001001001000000001111111111111110001111111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111111001111111111111111111111",
                  "1111111011011001111111111100001100110000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111111111000011111111111111111111111111111111111111001001001000000001111111111111110000111111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111111000111111111111111111111",
                  "1111111011011000000000000000111001100000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000000011000001111111111111111111111111111111111111001001001000000000000000000000010000011111100100100000000000000000000001001000000011110011011011000000111101101101100000001110010010011000000111100100100000000000000000000011111111111111111111",
                  "1111111011011111111111111111100011100000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000000011000000111111111111111111111111111111111111001001001000000000000000000000010000001111100100111111111111111111111111001000000011110011011011000000111101101101100000001110010010011000000111100100111111111111111110000000111111111111111111",
                  "1111111011011111111111111110000110000000000001110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111111011000000111111111111111111111111111111111111001001001000000001111111111110010000000111100100111111111111111111111111001000000011110011011011000000111101101101100000001110010010011000000111100100111111111111111111000000111111111111111111",
                  "1111111011011000000000000000011100000000000011110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000011011000000111111111111111111111111111111111111001001001000000000000000000010010000000111100100100000000000000000000001001000000011110011011011000000111101101101100000001110010010011000000111100100100000000000000000000000111111111111111111",
                  "1111111011011001111111111111110000000000000011110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000000011011000000111111111111111111111111111111111111001001001000000000000000000010010000000111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111110000000111111111111111111",
                  "1111111011011011111111111110000000000000000111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000001111111111011011000000111111111111111111111111111111111111001001001000000001111111110010010000000111100100100111111111111111111001001000000011110011011011000000111101101101100000001110010010011000000111100100100111111111111111000000111111111111111111",
                  "1111111011011011000000000000000000000000001111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000011011011000000111111111111111111111111111111111111001001001000000000000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000000011111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000011011011000000111111111111111111111111111111111111001001001000000000000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000000111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000000000000011011011000000111111111111111111111111111111111111001001001000000010000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000001111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011000000011011011000000111111111111111111111111111111111111001001001000000011000000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000000111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011100000011011011000000111111111111111111111111111111111111001001001000000011100000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000000011111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011110000011011011000000111111111111111111111111111111111111001001001000000011110000010010010000000111100100100100000000000000001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000111111111111111111",
                  "1111111011011011000000000000000011111111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111000011011011000000111111111111111111111111111111111111001001001000000011111000010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000000000000000000000000111111111111",
                  "1111111011011011000000011111111111111111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111110011011011000000111111111111111111111111111111111111001001001000000011111110010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111001000000100011111111111",
                  "1111111011011011000000011111111111111111111111110110110010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111110011011011000000111111111111111111111111111111111111001001001000000011111110010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100100000001111111001101101100001111111111",
                  "1111111011011011000000011111111111111111111111110110010010000000111111101101100100000001111011011001000000011111110110110010000000111001001101100000011111110010011011000000111111111111111111111111111111111111001001001000000011111110010010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100100110000001111111011001101100000111111111",
                  "1111111011011011000000011111111111111111111111110010010011000000111111001001101100000001111011011001000000011111110110110010000000111001101100100000011111110010010010000000111111111111111111111111111111111111001001101100000011111110110010010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100100110110000001111110011001001100000011111111",
                  "1111111011011011000000011111111111111111111111110010011011000000111111001001001100000001111011011001000000011111110110110010000000111101100100100000011111110110010010000000111111111111111111111111111111111111001101100100000011111100110110010000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111100110110010000001111110011001001000000011111111",
                  "1111111011011011000000011111111111111111111111110011001001100000111110011011001000000001111011011001000000011111110110110010000000111100100110110000011111100100110010000000111111111111111111111111111111111111101100100110000011111000100110110000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111110110010011000001111100110011011000000001111111",
                  "1111111011011011000000011111111111111111111111111011001001110000111000010011011000000001111011011001000000011111110110110010000000111100110110011000011110001100100110000000111111111111111111111111111111111111100100110010000011110001000100100000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111110010011001100001110001110010011000000001111111",
                  "1111111011011011000000011111111111111111111111111001100100111000000001100110011000000001111011011001000000011111110110110010000000111110010011001100000000011001100100000000111111111111111111111111111111111111100110011001100000000010001101100000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111110011001100110000000011100110110000000001111111",
                  "1111111011011011000000011111111111111111111111111001100110011110001111001100110000000001111011011001000000011111110110110010000000111110011001100111100011110011001100000000111111111111111111111111111111111111110010001000111100011100011001000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111001100110001111111110001100110000000011111111",
                  "1111111011011011000000011111111111111111111111111100110011000111111100011100100000000001111011011001000000011111110110110010000000111111001100110001111111000110011000000000111111111111111111111111111111111111110011001110001111110000110011000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111100100011000001111000011001100000000011111111",
                  "1111111011011011000000011111111111111111111111111110011001100000000000111001100000000011111011011001000000011111110110110010000000111111000110011100000000001100010000000000111111111111111111111111111111111111111001100011000000000001100110000000000111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111100110001110000000001110011000000000011111111",
                  "1111111011011011000000011111111111111111111111111110001100011100000111100011000000000011111011011001000000011111110110110010000000111111100011001111000001111000100000000000111111111111111111111111111111111111111100110001111000001110001100000000001111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111110011100111111111111000110000000000011111111",
                  "1111111011011011000000011111111111111111111111111111000110001111111110001110000000000011111011011001000000011111110110110010000000111111110001100011111111100011000000000001111111111111111111111111111111111111111110011100011111111000011000000000001111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111000110000111111100011100000000000111111111",
                  "1111111011011011000000011111111111111111111111111111100011100000000000011100000000000111111011011001000000011111110110110010000000111111111000111000000000000110000000000001111111111111111111111111111111111111111111000110000000000001110000000000001111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111100011100000000001111000000000000111111111",
                  "1111111011011011000000011111111111111111111111111111110001111000000011110000000000000111111011011001000000011111110110110010000000111111111100011111000001111100000000000011111111111111111111111111111111111111111111100011110000001111000000000000011111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111110000111111111111100000000000001111111111",
                  "1111111011011011000000011111111111111111111111111111111100001111111111000000000000001111111011011001000000011111110110110010000000111111111110000011111111100000000000000011111111111111111111111111111111111111111111110000111111111100000000000000111111100100100100000001111111001001001000000011110011011011000000111101101101100000001110010010011000000111111111111000000111111100000000000000001111111111",
                  "1111111000000000000000011111111111111111111111111111111110000000000000000000000000011111111000000000000000011111110000000000000000111111111111000000000000000000000000000111111111111111111111111111111111111111111111111000000000000000000000000000111111100000000000000001111111000000000000000011110000000000000000111100000000000000001110000000000000000111111111111100000000000000000000000000011111111111",
                  "1111111000000000000000011111111111111111111111111111111111000000000000000000000000011111111000000000000000011111110000000000000000111111111111100000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000001111111100000000000000001111111000000000000000011111000000000000000111100000000000000001110000000000000000111111111111110000000000000000000000000111111111111",
                  "1111111100000000000000011111111111111111111111111111111111100000000000000000000000111111111100000000000000011111111000000000000000111111111111110000000000000000000000011111111111111111111111111111111111111111111111111110000000000000000000000011111111110000000000000001111111110000000000000011111100000000000000111110000000000000001111100000000000000111111111111111100000000000000000000001111111111111",
                  "1111111110000000000000011111111111111111111111111111111111110000000000000000000011111111111110000000000000011111111100000000000000111111111111111100000000000000000000111111111111111111111111111111111111111111111111111111000000000000000000000111111111111000000000000001111111111000000000000011111110000000000000111111000000000000001111110000000000000111111111111111110000000000000000000011111111111111",
                  "1111111111000000000000011111111111111111111111111111111111111000000000000000000111111111111111000000000000011111111110000000000000111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000011111111111111100000000000001111111111100000000000011111111000000000000111111100000000000001111111000000000000111111111111111111000000000000000001111111111111111",
                  "1111111111100000000000011111111111111111111111111111111111111110000000000000011111111111111111100000000000011111111111000000000000111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111110000000000001111111111110000000000011111111100000000000111111110000000000001111111100000000000111111111111111111110000000000000111111111111111111",
                  "1111111111110000000000111111111111111111111111111111111111111111100000000011111111111111111111110000000000111111111111100000000000111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111100000000001111111111111000000000011111111110000000000111111111000000000011111111110000000000111111111111111111111111000001111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
    --The process involves the next state logic for the variables
    process(clock)
    begin 
        if clock'event and clock = '1' then
        --Producing the clock signal that will occur in the BallController module
            if ballMovementCounter = PRESCALER_BALL then
                ballMovement <= not ballMovement;
                ballMovementCounter <= 0;
            else 
                ballMovementCounter <= ballMovementCounter + 1;
            end if;
            --Button - paddle control
            if playing = '1' then
                if right = '1' and left = '0' then
                    paddleRight <= paddleRight + 1;
                    paddleLeft <= 0;
                elsif left = '1' and right = '0' then
                    paddleLeft <= paddleLeft + 1;
                    paddleRight <= 0;
                else 
                    paddleRight <= 0;
                    paddleLeft <= 0;
                end if;
                --Adjusting the position of the player's paddle according to the specified constant to avoid debouncing
                if paddleRight = (PRESCALER_PADDLE - 5000) and paddleCursor < TOT_H - paddleWidth then
                    paddleCursor <= paddleCursor + 1;
                elsif paddleLeft = (PRESCALER_PADDLE - 5000) and paddleCursor > FP_H + SP_H + BP_H + 1 then
                    paddleCursor <= paddleCursor - 1;
                end if;  
                --The basic A.I algorithm fot the computer to control a paddle, it follows the ball with a little pseudorandom error   
                if ballCursorX >= paddleAICursor + (ballCursorY mod (ballCursorX mod 5)) * ((ballCursorX) mod (ballCursorY mod 5)) + (paddleCursor * paddleAICursor) mod 5 then
                    paddleAIRight <= paddleAIRight + 1;
                    paddleAILeft <= 0;
                elsif ballCursorX <= paddleAICursor - (ballCursorY mod (ballCursorX mod 5)) * ((ballCursorX) mod (ballCursorY mod 5)) - (paddleCursor * paddleAICursor) mod 5 then 
                    paddleAILeft <= paddleAILeft + 1;
                    paddleAIRight <= 0;
                else 
                    paddleAILeft <= 0;
                    paddleAIRight <= 0;
                end if;
                --Adjusting the position of the computer's paddle according to the specified constant to avoid debouncing    
                if paddleAIRight = PRESCALER_PADDLE and paddleAICursor < TOT_H - PADDLE_WIDTH then
                    paddleAICursor <= paddleAICursor + 1;
                elsif paddleAILeft = PRESCALER_PADDLE and paddleAICursor > FP_H + SP_H + BP_H + 1 then
                    paddleAICursor <= paddleAICursor - 1;
                end if;                
            else --The initial positions of the paddles when the game stops
                paddleCursor <= FP_H + SP_H + BP_H + VIS_H / 2 - (PADDLE_WIDTH + 1) / 2;
                paddleAICursor <= FP_H + SP_H + BP_H + VIS_H / 2 - (PADDLE_WIDTH + 1) / 2;
            end if;
            --Register to update the values of the synchronization adn rgb signals
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
        end if;
    end process;
    --Difficulty selection with a multiplexer
    with difficultyControl select paddleWidth <= 
        PADDLE_WIDTH when "00",
        PADDLE_WIDTH_EASY when "01",
        PADDLE_WIDTH_HARD when "10",
        PADDLE_WIDTH when others;  
    --Cursor Position Selections
    result1Visible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 135) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 74) and
                      (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 150) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 150) and
                       result1(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 135))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 150)) 
                       = '0' and AIWins = '1';                  
    result2Visible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 135) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 74) and
                      (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 150) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 150) and
                      result2(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 135))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 150)) 
                      = '0' and playerWins = '1';
    messageVisible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 50) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 3) and
                      (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 200) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 200) and
                       message(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 50))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 200)) 
                       = '0' and newGame = '1';
    logoVisible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) + 45) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) + 210) and
                   (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 100) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 100) and
                    logo(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) + 45))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 100)) 
                    = '0' and newGame = '1';
    gameLabelVisible <= (vPosCurrent >= FP_V + SP_V + BP_V + (VIS_V / 2) - 138) and (vPosCurrent < FP_V + SP_V + BP_V + (VIS_V / 2) - 74) and
                        (hPosCurrent >= FP_H + SP_H + BP_H + (VIS_H / 2) - 200) and (hPosCurrent < FP_H + SP_H + BP_H + (VIS_H / 2) + 200) and
                        gameLabel(vPosCurrent - (FP_V + SP_V + BP_V + (VIS_V / 2) - 138))(hPosCurrent - (FP_H + SP_H + BP_H + (VIS_H / 2) - 200)) 
                        = '0' and AIWins = '0' and playerWins = '0' and newGame = '1';                                                                          
    paddleVisible <= ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 1) and (hPosCurrent > paddleCursor + 8) and (hPosCurrent < paddleCursor + paddleWidth - 8)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 1) and (hPosCurrent > paddleCursor + 7) and (hPosCurrent < paddleCursor + paddleWidth - 7)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 2) and (hPosCurrent > paddleCursor + 6) and (hPosCurrent < paddleCursor + paddleWidth - 6)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 3) and (hPosCurrent > paddleCursor + 5) and (hPosCurrent < paddleCursor + paddleWidth - 5)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 4) and (hPosCurrent > paddleCursor + 4) and (hPosCurrent < paddleCursor + paddleWidth - 4)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 5) and (hPosCurrent > paddleCursor + 3) and (hPosCurrent < paddleCursor + paddleWidth - 3)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 6) and (hPosCurrent > paddleCursor + 2) and (hPosCurrent < paddleCursor + paddleWidth - 2)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 7) and (hPosCurrent > paddleCursor + 1) and (hPosCurrent < paddleCursor + paddleWidth - 1)) or
                     (((vPosCurrent = TOT_V - PADDLE_HEIGHT + 8) or (vPosCurrent = TOT_V - PADDLE_HEIGHT + 9) or (vPosCurrent = TOT_V - PADDLE_HEIGHT + 10)) 
                     and (hPosCurrent > paddleCursor) and (hPosCurrent < paddleCursor + paddleWidth)) or
                     ((vPosCurrent = TOT_V - PADDLE_HEIGHT + 11) and (hPosCurrent > paddleCursor + 1) and (hPosCurrent < paddleCursor + paddleWidth - 1));
    ballVisible <= (((vPosCurrent = ballCursorY) or (vPosCurrent = ballCursorY + BALL_SIDE)) and (hPosCurrent > ballCursorX + 3) and (hPosCurrent <= ballCursorX + 7)) or
                   (((vPosCurrent = ballCursorY + 1) or (vPosCurrent = ballCursorY + BALL_SIDE - 1)) and (hPosCurrent > ballCursorX + 1) and (hPosCurrent <= ballCursorX + 9)) or
                   (((vPosCurrent = ballCursorY + 2) or (vPosCurrent = ballCursorY + BALL_SIDE - 2)
                   or (vPosCurrent = ballCursorY + 3) or (vPosCurrent = ballCursorY + BALL_SIDE - 3)) and (hPosCurrent > ballCursorX) and (hPosCurrent <= ballCursorX + 10)) or
                   ((vPosCurrent > ballCursorY + 2) and (vPosCurrent <= ballCursorY + 7) and (hPosCurrent >= ballCursorX) and (hPosCurrent <= ballCursorX + 11));
    paddleAIVisible <= ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 11) and (hPosCurrent > paddleAICursor + 8) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 8)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 10) and (hPosCurrent > paddleAICursor + 7) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 7)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 9) and (hPosCurrent > paddleAICursor + 6) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 6)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 8) and (hPosCurrent > paddleAICursor + 5) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 5)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 7) and (hPosCurrent > paddleAICursor + 4) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 4)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 6) and (hPosCurrent > paddleAICursor + 3) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 3)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 5) and (hPosCurrent > paddleAICursor + 2) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 2)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1 + 4) and (hPosCurrent > paddleAICursor + 1) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 1)) or
                       (((vPosCurrent = FP_V + SP_V + BP_V + 1 + 3) or (vPosCurrent = FP_V + SP_V + BP_V + 1 + 2) or (vPosCurrent = FP_V + SP_V + BP_V + 1 + 1)) 
                       and (hPosCurrent > paddleAICursor) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH)) or
                       ((vPosCurrent = FP_V + SP_V + BP_V + 1) and (hPosCurrent > paddleAICursor + 1) and (hPosCurrent < paddleAICursor + PADDLE_WIDTH - 1));                                          
    borderVisible <= (vPosCurrent = FP_V + SP_V + BP_V + (VIS_V / 2) and newGame = '0');
    --Scanning the Pixels
    hPosNext <= hPosCurrent + 1 when hPosCurrent < TOT_H else 1;
    vPosNext <= vPosCurrent + 1 when hPosCurrent = TOT_H and vPosCurrent < TOT_V else
                1 when hPosCurrent = TOT_H and vPosCurrent = TOT_V else vPosCurrent;
	--Color Selection with a multiplexer
    rgbNext <= "001011110001" when paddleVisible else
               "001110100010" when messageVisible else
               "001101111111" when ballVisible else                     
               "000000001111" when frameVisible or borderVisible else
               "011010010001" when paddleAIVisible else
               "100101000100" when result1Visible else
               "000010101110" when result2Visible else
               "001001101110" when gameLabelVisible else
               "000010101110" when logoVisible else
               "000000000000";    
    --Updating the signals that will go to the VGA port
    hSync <= '0' when (hPosCurrent > FP_H) and (hPosCurrent < FP_H + SP_H + 1) else '1';
    vSync <= '0' when (vPosCurrent > FP_V) and (vPosCurrent < FP_V + SP_V + 1) else '1';
    r <= rgbCurrent(11 downto 8);
    g <= rgbCurrent(7 downto 4);
    b <= rgbCurrent(3 downto 0);    
end Behavioral;
